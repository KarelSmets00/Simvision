*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.  
*/////////////////////////////////////////////////////////////////////
* Legal Notice:  
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice. 
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND" 
*////////////////////////////////////////////////////////////////////
*LMV7219 7nsec 2.7 to 5V Comparator with Rail-to-Rail Output
simulator lang = pspice

* PINOUT ORDER   +IN -IN VCC VSS OUT
.SUBCKT LMV7219   22  6   1   2  18
R1 1 3 10.0E6
V3 49 2 -1.2
V5 4 6 0.001
V4 1 42 0.6
Q1 47 47 42 Q1M
I3 47 2 40.0E-6
V15 48 2 -1.2
I2 1 2 2.1E-3
D1 50 46 D1M 
R3 5 46 3.5E6
R2 1 2 11.4E3
E6 43 0 30 0 1.0
E7 28 0 32 0 1.0
E8 8 0 26 0 1.0
G1 0 10 46 27 0.01
R6 10 0 100.0
R7 10 9 10.0
C5 9 0 62.0E-12
G2 0 11 10 0 -22.7E-3
R8 11 0 14.0E6
D5 12 11 DN4
D6 11 12 DN4
E1 12 0 13 0 1.0
R9 11 13 74.0
C6 13 0 0.05E-12
G3 0 14 13 0 0.01
R10 14 0 100.0
M1 18 14 1 1 WPM L=100U W=100U
M2 18 14 2 2 WNM L=100U W=100U
RO1 1 18 200.0E6
RO2 2 18 100.0E6
C1 14 0 10.0E-12
R14 46 24 1.0E9
R15 5 24 1.0E9
G6 0 26 24 0 5.6E-4
D8 34 1 D8M
V9 34 38 0.7
C2 14 18 1.0E-14
C3 18 0 1.0E-13
E2 16 0 14 0 1.0
RD3 16 0 1.0E18
E10 15 16 1 2 -0.7
R4 33 15 750.0
R16 26 25 1.0
L1 25 0 3.2E-8
E3 5 27 39 0 1.0
I1 0 37 1.0E-3
G7 0 32 2 0 6.0E-5
G8 0 30 1 0 6.0E-5
R24 30 29 1.0
L2 29 0 1.6E-7
R25 32 31 1.0
L3 31 0 1.6E-7
V13 41 37 -0.71465
D15 40 36 D8M 
V12 13 36 0.7
E4 39 0 0 33 1.0E6
R29 33 43 1.0
R30 33 28 1.0
R31 33 8 1.0
R32 39 33 1.0
E5 38 13 41 0 1.0
E9 40 2 41 0 1.0
D10 37 0 D8M
D2 52 5 D1M
Q3 3 47 42 QAM 10
R19 3 44 1.0E3
R20 3 45 999.0
R22 46 48 1.0E3
R23 5 49 999.0
Q4 50 4 44 Q4M
Q5 52 22 45 Q5M
RD1 27 0 1.0E18
RD2 41 0 1.0E18
.MODEL D8M D IS=1.0E-15
.MODEL DN4 D BV=100.0 CJO=4.0E-12 IS=7.0E-9
+ M=0.45 N=2 RS=0.8 TT=6.0E-9 VJ=0.6
.MODEL D1M D BV=5.33E+1 CJO=2.0E-14
+ IBV=5.0E-8 IS=4.69E-16 M=0.333 N=1.95
+ RS=2.18E-1 TT=2.9E-9 VJ=0.75
.MODEL Q1M PNP BF=200.0
.MODEL QAM PNP BF=100.0
.MODEL Q4M PNP BF=200.0
.MODEL Q5M PNP BF=250.0
.MODEL WNM NMOS LEVEL=1 KP=0.015 RD=32.0 RS=1.0
+ VTO=1.0 IS=1.0E-14 FC=0.5 MJ=0.5 MJSW=0.5 PB=0.8
+ PHI=0.6 TOX=1.0E-7 UO=600.0 TPG=1 AF=1
.MODEL WPM PMOS LEVEL=1 KP=0.015 RD=32.0 RS=1.0
+ VTO=-1.0 IS=1.0E-14 FC=0.5 MJ=0.5 MJSW=0.5 PB=0.8
+ PHI=0.6 TOX=1.0E-7 UO=600.0 TPG=1 AF=1
.ENDS

