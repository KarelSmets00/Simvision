`timescale 1ns/1ps

module Counter (
	input wire clk,
	input wire nrst,
	input wire enable,
	output reg [7:0] value
	);


	

endmodule
