`timescale 1ns/1ps


module toplevel ();

	ANALOG_NETWORK analog_network_inst (
	);

endmodule
