simulator lang = spice
.param D=0.5
.param P=0.0126m

.SUBCKT ANALOG_NETWORK 
.option post=1

.param Von=3.3

.param k12=0.605 k23=0.082746 k34=0.62499 k13=0.065501 k14=0.051516 k24=0.064887
.param LL1=2.6567e-05 LL2=0.00044945 LL3=0.00063979 LL4=3.6751e-05
.param RR1=0.11647 RR2=0.56704 RR3=0.75095 RR4=0.15326
.param CC1=3.8139e-07 CC2=2.2543e-08 CC3=1.5837e-08 CC4=2.757e-07

.param Rm=100

.include DI_BAV5004LP.spi

XX1 3v3 0 N008 N011 0 12v 0 N010 N016 N013 N019 h_bridge
V1 3v3 0 3.3
V2 12v 0 12 Rser=0
XX2 N008 N011 N013 N019 pwm_sourcev2
XX4 N007 N017 VDC 0 full_bridge_rect
C1 VDC 0 100u
R1 VDC 0 80
L1 N009 N016 LL1
L2 N014 N002 LL2
L3 N006 N015 LL3
L4 N017 N004 LL4
C2 N005 N014 CC2
C3 N003 N015 CC3
R9 N005 N002 RR2
R10 N006 N003 RR3
C4 N007 N017 CC4
C5 N010 N001 CC1
R11 N001 N009 RR1
R12 N007 N004 RR4
R13 N002 N001 1G
R14 N003 N005 1G
R15 N004 N006 1G
V3 5Vrx 0 5V
D5 N007 ENV DI_BAV5004LP
D6 N017 ENV DI_BAV5004LP
C6 ENV 0 0.62u
R16 ENV 0 1k
C7 ENV MOD 1u
R17 MOD 0 1.5k


K12 L1 L2 k12
K23 L2 L3 k23
K34 L3 L4 k34
K14 L1 L4 k14
K13 L1 L3 k13
K24 L2 L4 k24

* block symbol definitions

.subckt h_bridge Vlog SD G1 G2 LGND Vcc COMM ACL ACN G3 G4
XU1 Vlog G1 SD G3 LGND N001 N003 ACL Vcc COMM N005 IR2110
XU2 Vcc N001 ACL irfs_sl7440pbf
XU3 ACL N005 COMM irfs_sl7440pbf
XU4 Vcc N002 ACN irfs_sl7440pbf
XU5 ACN N006 COMM irfs_sl7440pbf
XU6 Vlog G2 SD G4 LGND N002 N004 ACN Vcc COMM N006 IR2110
C1 N003 ACL 500n
D5 Vcc N003 DI_BAV5004LP
C2 COMM Vcc 10n
C3 N004 ACN 500n
D6 Vcc N004 DI_BAV5004LP
C4 Vcc COMM 10n
C5 Vlog LGND 10n
C6 Vlog LGND 10n
.include DI_BAV5004LP.spi
.include IR2110.spi
.include irfs_sl7440pbf.spi
.ENDS

.subckt pwm_sourcev2 G1 G2 G3 G4
V1 G1 0 PULSE(0 Von 0 0.1n 0.1n P*D P*2)
V2 G2 0 PULSE(0 Von P 0.1n 0.1n P*D P*2)
E1 G3 N001 G1 0 -1
E2 G4 N002 G2 0 -1
V3 N001 0 Von
V4 N002 0 Von
.ENDS

.subckt full_bridge_rect ACL ACN V+ V-
D1 ACN V+ d1n5408
D2 ACL V+ d1n5408
D3 V- ACN d1n5408
D4 V- ACL d1n5408
.include 1N5408.spi
.ENDS



* PARAMETERS\nberekend op resonantiefrequentie = 50kHz\noptimale overdracht op freq = 39267.2 Hz\nwss best om H-brug aan te sturen op die frequentie. \n \n.param k12=0.62499 k23=0.10311 k34=0.62499 k13=0.081644 k14=0.064839 k24=0.081644\n.param L1=3.6751e-05 L2=0.00063979 L3=0.00063979 L4=3.6751e-05\n.param R1=0.15326 R2=0.75095 R3=0.75095 R4=0.15326\n.param C1=2.757e-07 C2=1.5837e-08 C3=1.5837e-08 C4=2.757e-07


.ENDS

simulator lang = spectre
