*******************************************************************
* Model name       : BAT48
* Description      : Small Signal Schottky Diode
* Package type     : DO35
*******************************************************************
.MODEL BAT48 D IS=263.91E-9 N=1.0966 RS=.4109 IKF=29.589E-3
+ EG=.69 XTI=2 CJO=29.800E-12 M=.50094 VJ=.41054 ISR=90.294E-9
+ FC=0.5 NR=4.9949 TT=0
