simulator lang = spice

.SUBCKT ANALOG_NETWORK 
.option post=1

.param Rled=28.8
.param Rcirc=15

.param k12=0.62499 k23=0.10311 k34=0.62499 k13=0.081644 k14=0.064839 k24=0.081644
.param LL1=3.6751e-05 LL2=0.00063979 LL3=0.00063979 LL4=3.6751e-05
.param RR1=0.15326 RR2=0.75095 RR3=0.75095 RR4=0.15326
.param CC1=2.757e-07 CC2=1.5837e-08 CC3=1.5837e-08 CC4=2.757e-07

.param P=0.01m
.param D=0.5
.param Von=3.3

.param Rm=100

.include OPA2344.spi
.include LM7812.spi
.include DI_10A01.spi


RLED_WALL +12V 0 Rled
C2 +12V 0 0.1u
C3 Vdc 0 4.7u
RCirc 5Vrx 0 Rcirc
XU2 Vdc 0 +12V LM7812
XX1 N005 N008 N006 0 full_bridge_rect
RNano 5Vrx 0 250
RLCD 5Vrx 0 125
XX2 5Vtx 0 N003 N007 0 Vbatt N013 N004 N011 N009 N012 h_bridge
XU3 N015 Ref 5Vtx 0 Ref OPA2344
R3 5Vtx N015 20k
R4 N015 0 5k
XX4 Vadc Vbatt 0 5Vtx Ref 0 dc_voltage
XX5 N013 0 Iadc 5Vtx Ref 0 dc_current
V2 Vbatt 0 11
XX6 Vbatt 5Vtx 0 dc_supply5v0
XX7 N004 N010 N005 N008 link_optimized
XX8 N003 N007 N009 N012 pwm_sourcev2 params: D=0.5,P=0.0127m,Von=5
XX3 N010 N011 Ref 0 5Vtx +Iac -Iac current_sensorv3
XX9 Vdc 5Vrx 0 dc_supply5v0
D1 N006 Vdc DI_10A01
C1 Vdc 0 100u
XX11 5Vrx 0 N006 Freq\ Freq freq_detect


.SUBCKT full_bridge_rect ACL ACN V+ V-
D1 ACN V+ DI_10A01
D2 ACL V+ DI_10A01
D3 V- ACN DI_10A01
D4 V- ACL DI_10A01
.include DI_10A01.spi
.ENDS

.SUBCKT h_bridge Vlog SD G1 G2 LGND Vcc COMM ACL ACN G3 G4
XU1 Vlog G1 SD G3 LGND N001 N003 ACL Vcc COMM N005 IR2110
XU2 Vcc N001 ACL irfs_sl7440pbf
XU3 ACL N005 COMM irfs_sl7440pbf
XU4 Vcc N002 ACN irfs_sl7440pbf
XU5 ACN N006 COMM irfs_sl7440pbf
XU6 Vlog G2 SD G4 LGND N002 N004 ACN Vcc COMM N006 IR2110
C1 N003 ACL 500n
D5 Vcc N003 DI_BAV5004LP
C2 COMM Vcc 10n
C3 N004 ACN 500n
D6 Vcc N004 DI_BAV5004LP
C4 Vcc COMM 10n
C5 Vlog LGND 10n
C6 Vlog LGND 10n
.include DI_BAV5004LP.spi
.include IR2110.spi
.include irfs_sl7440pbf.spi
.ENDS

.SUBCKT dc_voltage ADC Vin COMM Vdd INmax Agnd
R1 Vin N001 200k
R2 N001 COMM 10k
R3 N003 N002 100
XU1 N001 N002 Vdd COMM N002 OPA2344
D1 N004 INmax BAT48
D2 Agnd N004 BAT48
R4 ADC N003 100
.include OPA2344.spi
.include ST_BAT48.spi
.ENDS

.SUBCKT dc_current LOAD COMM ADC Vdd INmax Agnd
Rshunt LOAD COMM 10m
XU1 LOAD COMM Vdd COMM N001 INA180A1
R1 N002 N001 100
D1 N002 INmax BAT48
D2 Agnd N002 BAT48
R2 ADC N002 100
.include ina180a1.spi
.include ST_BAT48.spi
.ENDS

.SUBCKT dc_supply5v0 Vin 5V0 COMM
XU1 Vin N001 COMM N002 COMM COMM COMM COMM COMM COMM COMM COMM COMM COMM COMM COMM LM2575_TRANS
C1 Vin COMM 100u
L1 N001 5V0 330u
C2 5V0 COMM 330u
R1 5V0 N002 31k
R2 N002 COMM 10k
D1 COMM N001 D1n5819
.include LM2575_TRANS.spi
.include 1N5819.spi
.ENDS

.SUBCKT link_optimized IN1 IN2 OUT1 OUT2
L1 N007 IN2 LL1
L2 N008 N002 LL2
L3 N006 N009 LL3
L4 OUT2 N004 LL4
C1 N005 N008 CC2
C2 N003 N009 CC3
R1 N005 N002 RR2
R2 N006 N003 RR3
C3 OUT1 OUT2 CC4
C4 N001 IN1 CC1
R3 N001 N007 RR1
R4 OUT1 N004 RR4
R6 N002 N001 1G
R7 N003 N005 1G
R8 N004 N006 1G
K12 L1 L2 k12
K23 L2 L3 k23
K34 L3 L4 k34
K14 L1 L4 k14
K13 L1 L3 k13
K24 L2 L4 k24
.ENDS

.SUBCKT pwm_sourcev2 G1 G2 G3 G4
V1 G1 0 PULSE(0 {Von} 0 0 0 {P*D} {P*2})
V2 G2 0 PULSE(0 {Von} {P} 0 0 {P*D} {P*2})
E1 G3 N001 G1 0 -1
E2 G4 N002 G2 0 -1
V3 N001 0 {Von}
V4 N002 0 {Von}
.ENDS

.SUBCKT current_sensorv3 Cin Cout INmax Agnd Vcc ADC+ ADC-
F1 N002 N001 V1 1/Rm
R1 N001 Vcm 1Meg
R2 Vcm N002 1Meg
R3 Vcm Agnd 12k
R4 Vcc Vcm 100k
R5 N001 N002 10
V1 Cin Cout 0
R6 ADC+ N001 100
R7 ADC- N002 100
D1 ADC+ INmax BAT48
D2 ADC- INmax BAT48
D3 Agnd ADC+ BAT48
D4 Agnd ADC- BAT48
.include ST_BAT48.spi
.ENDS

.SUBCKT freq_detect Vcc COMM In+ Out\ Out
R1 In+ N001 10k
R2 N001 COMM 1k
XU1 N001 COMM Vcc COMM Out\ LMV7219
XU2 Out Out\ Out\ Vcc COMM SN74HC00
.include LMV7219.spi
.include SN74HC00.spi
.ENDS


.ENDS

simulator lang = spectre
