simulator lang = spice

.param freq = 50k

.SUBCKT ANALOG_NETWORK 
.option post=1

.include "SmallSignalDiode.spi"

VSS vss 0 0
Vpulse n1 vss SIN(0 12 freq)

D1 n1 n2 SmallSignalDiode
R1 n2 vss 100

Vfreq param_freq vss freq

.ENDS

simulator lang = spectre
